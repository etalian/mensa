VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_bfloat16
  CLASS BLOCK ;
  FOREIGN wrapped_bfloat16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.410 296.000 23.970 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.420 300.000 1.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.980 300.000 64.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 69.100 300.000 70.300 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 75.900 300.000 77.100 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 82.020 300.000 83.220 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.140 300.000 89.340 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.260 300.000 95.460 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.060 300.000 102.260 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.180 300.000 108.380 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 113.300 300.000 114.500 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.420 300.000 120.620 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 6.540 300.000 7.740 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 126.220 300.000 127.420 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 132.340 300.000 133.540 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.460 300.000 139.660 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.580 300.000 145.780 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.380 300.000 152.580 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.500 300.000 158.700 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.620 300.000 164.820 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.740 300.000 170.940 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.540 300.000 177.740 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.660 300.000 183.860 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 12.660 300.000 13.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.780 300.000 189.980 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 194.900 300.000 196.100 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.700 300.000 202.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.820 300.000 209.020 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.940 300.000 215.140 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.060 300.000 221.260 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 226.860 300.000 228.060 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.980 300.000 234.180 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.780 300.000 19.980 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.580 300.000 26.780 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.700 300.000 32.900 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.820 300.000 39.020 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 43.940 300.000 45.140 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.740 300.000 51.940 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 56.860 300.000 58.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 67.060 300.000 68.260 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.180 300.000 74.380 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.980 300.000 81.180 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.100 300.000 87.300 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.220 300.000 93.420 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 98.340 300.000 99.540 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.140 300.000 106.340 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.260 300.000 112.460 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.380 300.000 118.580 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.500 300.000 124.700 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.620 300.000 11.820 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.300 300.000 131.500 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.420 300.000 137.620 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.540 300.000 143.740 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.660 300.000 149.860 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.460 300.000 156.660 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.580 300.000 162.780 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.700 300.000 168.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 173.820 300.000 175.020 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.620 300.000 181.820 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.740 300.000 187.940 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.740 300.000 17.940 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.860 300.000 194.060 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.980 300.000 200.180 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.780 300.000 206.980 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.900 300.000 213.100 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 218.020 300.000 219.220 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.140 300.000 225.340 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 230.940 300.000 232.140 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.060 300.000 238.260 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 22.860 300.000 24.060 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.660 300.000 30.860 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.780 300.000 36.980 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 41.900 300.000 43.100 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 48.020 300.000 49.220 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.820 300.000 56.020 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.940 300.000 62.140 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.460 300.000 3.660 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.140 300.000 72.340 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 77.940 300.000 79.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.060 300.000 85.260 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 90.180 300.000 91.380 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.300 300.000 97.500 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.100 300.000 104.300 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 109.220 300.000 110.420 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.340 300.000 116.540 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 121.460 300.000 122.660 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.580 300.000 9.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 128.260 300.000 129.460 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 134.380 300.000 135.580 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 140.500 300.000 141.700 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.620 300.000 147.820 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 153.420 300.000 154.620 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.540 300.000 160.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.660 300.000 166.860 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.780 300.000 172.980 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 178.580 300.000 179.780 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 184.700 300.000 185.900 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 14.700 300.000 15.900 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.820 300.000 192.020 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 196.940 300.000 198.140 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.740 300.000 204.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.860 300.000 211.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.980 300.000 217.180 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 222.100 300.000 223.300 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.900 300.000 230.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.020 300.000 236.220 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.820 300.000 22.020 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.620 300.000 28.820 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.740 300.000 34.940 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.860 300.000 41.060 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 45.980 300.000 47.180 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.780 300.000 53.980 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 58.900 300.000 60.100 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.930 0.000 6.490 4.000 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 256.100 300.000 257.300 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.100 4.000 121.300 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.750 0.000 106.310 4.000 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.810 296.000 134.370 300.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.010 0.000 143.570 4.000 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 296.000 150.010 300.000 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.550 296.000 166.110 300.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.300 300.000 267.500 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 0.000 181.290 4.000 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.420 300.000 273.620 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 241.140 300.000 242.340 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.580 4.000 213.780 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.220 300.000 280.420 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.930 296.000 213.490 300.000 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 283.300 300.000 284.500 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.340 300.000 286.540 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.570 0.000 206.130 4.000 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.990 0.000 218.550 4.000 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.820 4.000 260.020 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.290 0.000 243.850 4.000 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.130 0.000 268.690 4.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 243.180 300.000 244.380 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.500 300.000 294.700 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.540 300.000 296.740 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.620 4.000 28.820 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.190 0.000 43.750 4.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 0.000 68.590 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.740 4.000 51.940 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.860 4.000 75.060 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.420 4.000 86.620 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 0.000 93.890 4.000 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.180 4.000 6.380 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.140 300.000 259.340 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.180 300.000 261.380 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.660 4.000 132.860 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.590 0.000 131.150 4.000 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 262.220 300.000 263.420 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 264.260 300.000 265.460 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.340 4.000 167.540 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.340 300.000 269.540 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 270.380 300.000 271.580 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.020 4.000 202.220 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.140 4.000 225.340 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 296.000 181.750 300.000 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 0.000 193.710 4.000 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 296.000 229.130 300.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.700 4.000 236.900 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.380 300.000 288.580 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.590 296.000 292.150 300.000 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 0.000 231.430 4.000 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.380 4.000 271.580 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.460 300.000 292.660 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 296.000 55.250 300.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.940 4.000 283.140 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.500 4.000 294.700 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.770 0.000 31.330 4.000 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 0.000 56.170 4.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.180 4.000 40.380 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.790 296.000 71.350 300.000 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.430 296.000 86.990 300.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 0.000 81.470 4.000 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.100 300.000 240.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.170 296.000 118.730 300.000 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.170 0.000 118.730 4.000 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.220 4.000 144.420 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.890 0.000 156.450 4.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.780 4.000 155.980 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 0.000 168.870 4.000 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.900 4.000 179.100 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.460 4.000 190.660 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.460 300.000 275.660 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.050 296.000 39.610 300.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.180 300.000 278.380 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 296.000 197.390 300.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.260 300.000 282.460 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.210 296.000 244.770 300.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.310 296.000 260.870 300.000 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 296.000 276.510 300.000 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.260 4.000 248.460 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 0.000 256.270 4.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 0.000 281.110 4.000 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.060 4.000 17.260 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.970 0.000 293.530 4.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.580 300.000 298.780 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 245.220 300.000 246.420 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.260 300.000 248.460 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 249.300 300.000 250.500 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.070 296.000 102.630 300.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.020 300.000 253.220 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.060 300.000 255.260 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.770 296.000 8.330 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 5.520 10.640 294.400 288.560 ;
      LAYER met2 ;
        RECT 7.000 295.720 7.490 296.210 ;
        RECT 8.610 295.720 23.130 296.210 ;
        RECT 24.250 295.720 38.770 296.210 ;
        RECT 39.890 295.720 54.410 296.210 ;
        RECT 55.530 295.720 70.510 296.210 ;
        RECT 71.630 295.720 86.150 296.210 ;
        RECT 87.270 295.720 101.790 296.210 ;
        RECT 102.910 295.720 117.890 296.210 ;
        RECT 119.010 295.720 133.530 296.210 ;
        RECT 134.650 295.720 149.170 296.210 ;
        RECT 150.290 295.720 165.270 296.210 ;
        RECT 166.390 295.720 180.910 296.210 ;
        RECT 182.030 295.720 196.550 296.210 ;
        RECT 197.670 295.720 212.650 296.210 ;
        RECT 213.770 295.720 228.290 296.210 ;
        RECT 229.410 295.720 243.930 296.210 ;
        RECT 245.050 295.720 260.030 296.210 ;
        RECT 261.150 295.720 275.670 296.210 ;
        RECT 276.790 295.720 291.310 296.210 ;
        RECT 292.430 295.720 292.920 296.210 ;
        RECT 7.000 4.280 292.920 295.720 ;
        RECT 7.000 2.875 18.070 4.280 ;
        RECT 19.190 2.875 30.490 4.280 ;
        RECT 31.610 2.875 42.910 4.280 ;
        RECT 44.030 2.875 55.330 4.280 ;
        RECT 56.450 2.875 67.750 4.280 ;
        RECT 68.870 2.875 80.630 4.280 ;
        RECT 81.750 2.875 93.050 4.280 ;
        RECT 94.170 2.875 105.470 4.280 ;
        RECT 106.590 2.875 117.890 4.280 ;
        RECT 119.010 2.875 130.310 4.280 ;
        RECT 131.430 2.875 142.730 4.280 ;
        RECT 143.850 2.875 155.610 4.280 ;
        RECT 156.730 2.875 168.030 4.280 ;
        RECT 169.150 2.875 180.450 4.280 ;
        RECT 181.570 2.875 192.870 4.280 ;
        RECT 193.990 2.875 205.290 4.280 ;
        RECT 206.410 2.875 217.710 4.280 ;
        RECT 218.830 2.875 230.590 4.280 ;
        RECT 231.710 2.875 243.010 4.280 ;
        RECT 244.130 2.875 255.430 4.280 ;
        RECT 256.550 2.875 267.850 4.280 ;
        RECT 268.970 2.875 280.270 4.280 ;
        RECT 281.390 2.875 292.690 4.280 ;
      LAYER met3 ;
        RECT 4.400 293.100 295.600 294.265 ;
        RECT 4.000 293.060 296.000 293.100 ;
        RECT 4.000 291.060 295.600 293.060 ;
        RECT 4.000 291.020 296.000 291.060 ;
        RECT 4.000 289.020 295.600 291.020 ;
        RECT 4.000 288.980 296.000 289.020 ;
        RECT 4.000 286.980 295.600 288.980 ;
        RECT 4.000 286.940 296.000 286.980 ;
        RECT 4.000 284.940 295.600 286.940 ;
        RECT 4.000 284.900 296.000 284.940 ;
        RECT 4.000 283.540 295.600 284.900 ;
        RECT 4.400 282.900 295.600 283.540 ;
        RECT 4.400 282.860 296.000 282.900 ;
        RECT 4.400 281.540 295.600 282.860 ;
        RECT 4.000 280.860 295.600 281.540 ;
        RECT 4.000 280.820 296.000 280.860 ;
        RECT 4.000 278.820 295.600 280.820 ;
        RECT 4.000 278.780 296.000 278.820 ;
        RECT 4.000 276.780 295.600 278.780 ;
        RECT 4.000 276.060 296.000 276.780 ;
        RECT 4.000 274.060 295.600 276.060 ;
        RECT 4.000 274.020 296.000 274.060 ;
        RECT 4.000 272.020 295.600 274.020 ;
        RECT 4.000 271.980 296.000 272.020 ;
        RECT 4.400 269.980 295.600 271.980 ;
        RECT 4.000 269.940 296.000 269.980 ;
        RECT 4.000 267.940 295.600 269.940 ;
        RECT 4.000 267.900 296.000 267.940 ;
        RECT 4.000 265.900 295.600 267.900 ;
        RECT 4.000 265.860 296.000 265.900 ;
        RECT 4.000 263.860 295.600 265.860 ;
        RECT 4.000 263.820 296.000 263.860 ;
        RECT 4.000 261.820 295.600 263.820 ;
        RECT 4.000 261.780 296.000 261.820 ;
        RECT 4.000 260.420 295.600 261.780 ;
        RECT 4.400 259.780 295.600 260.420 ;
        RECT 4.400 259.740 296.000 259.780 ;
        RECT 4.400 258.420 295.600 259.740 ;
        RECT 4.000 257.740 295.600 258.420 ;
        RECT 4.000 257.700 296.000 257.740 ;
        RECT 4.000 255.700 295.600 257.700 ;
        RECT 4.000 255.660 296.000 255.700 ;
        RECT 4.000 253.660 295.600 255.660 ;
        RECT 4.000 253.620 296.000 253.660 ;
        RECT 4.000 251.620 295.600 253.620 ;
        RECT 4.000 250.900 296.000 251.620 ;
        RECT 4.000 248.900 295.600 250.900 ;
        RECT 4.000 248.860 296.000 248.900 ;
        RECT 4.400 246.860 295.600 248.860 ;
        RECT 4.000 246.820 296.000 246.860 ;
        RECT 4.000 244.820 295.600 246.820 ;
        RECT 4.000 244.780 296.000 244.820 ;
        RECT 4.000 242.780 295.600 244.780 ;
        RECT 4.000 242.740 296.000 242.780 ;
        RECT 4.000 240.740 295.600 242.740 ;
        RECT 4.000 240.700 296.000 240.740 ;
        RECT 4.000 238.700 295.600 240.700 ;
        RECT 4.000 238.660 296.000 238.700 ;
        RECT 4.000 237.300 295.600 238.660 ;
        RECT 4.400 236.660 295.600 237.300 ;
        RECT 4.400 236.620 296.000 236.660 ;
        RECT 4.400 235.300 295.600 236.620 ;
        RECT 4.000 234.620 295.600 235.300 ;
        RECT 4.000 234.580 296.000 234.620 ;
        RECT 4.000 232.580 295.600 234.580 ;
        RECT 4.000 232.540 296.000 232.580 ;
        RECT 4.000 230.540 295.600 232.540 ;
        RECT 4.000 230.500 296.000 230.540 ;
        RECT 4.000 228.500 295.600 230.500 ;
        RECT 4.000 228.460 296.000 228.500 ;
        RECT 4.000 226.460 295.600 228.460 ;
        RECT 4.000 225.740 296.000 226.460 ;
        RECT 4.400 223.740 295.600 225.740 ;
        RECT 4.000 223.700 296.000 223.740 ;
        RECT 4.000 221.700 295.600 223.700 ;
        RECT 4.000 221.660 296.000 221.700 ;
        RECT 4.000 219.660 295.600 221.660 ;
        RECT 4.000 219.620 296.000 219.660 ;
        RECT 4.000 217.620 295.600 219.620 ;
        RECT 4.000 217.580 296.000 217.620 ;
        RECT 4.000 215.580 295.600 217.580 ;
        RECT 4.000 215.540 296.000 215.580 ;
        RECT 4.000 214.180 295.600 215.540 ;
        RECT 4.400 213.540 295.600 214.180 ;
        RECT 4.400 213.500 296.000 213.540 ;
        RECT 4.400 212.180 295.600 213.500 ;
        RECT 4.000 211.500 295.600 212.180 ;
        RECT 4.000 211.460 296.000 211.500 ;
        RECT 4.000 209.460 295.600 211.460 ;
        RECT 4.000 209.420 296.000 209.460 ;
        RECT 4.000 207.420 295.600 209.420 ;
        RECT 4.000 207.380 296.000 207.420 ;
        RECT 4.000 205.380 295.600 207.380 ;
        RECT 4.000 205.340 296.000 205.380 ;
        RECT 4.000 203.340 295.600 205.340 ;
        RECT 4.000 203.300 296.000 203.340 ;
        RECT 4.000 202.620 295.600 203.300 ;
        RECT 4.400 201.300 295.600 202.620 ;
        RECT 4.400 200.620 296.000 201.300 ;
        RECT 4.000 200.580 296.000 200.620 ;
        RECT 4.000 198.580 295.600 200.580 ;
        RECT 4.000 198.540 296.000 198.580 ;
        RECT 4.000 196.540 295.600 198.540 ;
        RECT 4.000 196.500 296.000 196.540 ;
        RECT 4.000 194.500 295.600 196.500 ;
        RECT 4.000 194.460 296.000 194.500 ;
        RECT 4.000 192.460 295.600 194.460 ;
        RECT 4.000 192.420 296.000 192.460 ;
        RECT 4.000 191.060 295.600 192.420 ;
        RECT 4.400 190.420 295.600 191.060 ;
        RECT 4.400 190.380 296.000 190.420 ;
        RECT 4.400 189.060 295.600 190.380 ;
        RECT 4.000 188.380 295.600 189.060 ;
        RECT 4.000 188.340 296.000 188.380 ;
        RECT 4.000 186.340 295.600 188.340 ;
        RECT 4.000 186.300 296.000 186.340 ;
        RECT 4.000 184.300 295.600 186.300 ;
        RECT 4.000 184.260 296.000 184.300 ;
        RECT 4.000 182.260 295.600 184.260 ;
        RECT 4.000 182.220 296.000 182.260 ;
        RECT 4.000 180.220 295.600 182.220 ;
        RECT 4.000 180.180 296.000 180.220 ;
        RECT 4.000 179.500 295.600 180.180 ;
        RECT 4.400 178.180 295.600 179.500 ;
        RECT 4.400 178.140 296.000 178.180 ;
        RECT 4.400 177.500 295.600 178.140 ;
        RECT 4.000 176.140 295.600 177.500 ;
        RECT 4.000 175.420 296.000 176.140 ;
        RECT 4.000 173.420 295.600 175.420 ;
        RECT 4.000 173.380 296.000 173.420 ;
        RECT 4.000 171.380 295.600 173.380 ;
        RECT 4.000 171.340 296.000 171.380 ;
        RECT 4.000 169.340 295.600 171.340 ;
        RECT 4.000 169.300 296.000 169.340 ;
        RECT 4.000 167.940 295.600 169.300 ;
        RECT 4.400 167.300 295.600 167.940 ;
        RECT 4.400 167.260 296.000 167.300 ;
        RECT 4.400 165.940 295.600 167.260 ;
        RECT 4.000 165.260 295.600 165.940 ;
        RECT 4.000 165.220 296.000 165.260 ;
        RECT 4.000 163.220 295.600 165.220 ;
        RECT 4.000 163.180 296.000 163.220 ;
        RECT 4.000 161.180 295.600 163.180 ;
        RECT 4.000 161.140 296.000 161.180 ;
        RECT 4.000 159.140 295.600 161.140 ;
        RECT 4.000 159.100 296.000 159.140 ;
        RECT 4.000 157.100 295.600 159.100 ;
        RECT 4.000 157.060 296.000 157.100 ;
        RECT 4.000 156.380 295.600 157.060 ;
        RECT 4.400 155.060 295.600 156.380 ;
        RECT 4.400 155.020 296.000 155.060 ;
        RECT 4.400 154.380 295.600 155.020 ;
        RECT 4.000 153.020 295.600 154.380 ;
        RECT 4.000 152.980 296.000 153.020 ;
        RECT 4.000 150.980 295.600 152.980 ;
        RECT 4.000 150.260 296.000 150.980 ;
        RECT 4.000 148.260 295.600 150.260 ;
        RECT 4.000 148.220 296.000 148.260 ;
        RECT 4.000 146.220 295.600 148.220 ;
        RECT 4.000 146.180 296.000 146.220 ;
        RECT 4.000 144.820 295.600 146.180 ;
        RECT 4.400 144.180 295.600 144.820 ;
        RECT 4.400 144.140 296.000 144.180 ;
        RECT 4.400 142.820 295.600 144.140 ;
        RECT 4.000 142.140 295.600 142.820 ;
        RECT 4.000 142.100 296.000 142.140 ;
        RECT 4.000 140.100 295.600 142.100 ;
        RECT 4.000 140.060 296.000 140.100 ;
        RECT 4.000 138.060 295.600 140.060 ;
        RECT 4.000 138.020 296.000 138.060 ;
        RECT 4.000 136.020 295.600 138.020 ;
        RECT 4.000 135.980 296.000 136.020 ;
        RECT 4.000 133.980 295.600 135.980 ;
        RECT 4.000 133.940 296.000 133.980 ;
        RECT 4.000 133.260 295.600 133.940 ;
        RECT 4.400 131.940 295.600 133.260 ;
        RECT 4.400 131.900 296.000 131.940 ;
        RECT 4.400 131.260 295.600 131.900 ;
        RECT 4.000 129.900 295.600 131.260 ;
        RECT 4.000 129.860 296.000 129.900 ;
        RECT 4.000 127.860 295.600 129.860 ;
        RECT 4.000 127.820 296.000 127.860 ;
        RECT 4.000 125.820 295.600 127.820 ;
        RECT 4.000 125.100 296.000 125.820 ;
        RECT 4.000 123.100 295.600 125.100 ;
        RECT 4.000 123.060 296.000 123.100 ;
        RECT 4.000 121.700 295.600 123.060 ;
        RECT 4.400 121.060 295.600 121.700 ;
        RECT 4.400 121.020 296.000 121.060 ;
        RECT 4.400 119.700 295.600 121.020 ;
        RECT 4.000 119.020 295.600 119.700 ;
        RECT 4.000 118.980 296.000 119.020 ;
        RECT 4.000 116.980 295.600 118.980 ;
        RECT 4.000 116.940 296.000 116.980 ;
        RECT 4.000 114.940 295.600 116.940 ;
        RECT 4.000 114.900 296.000 114.940 ;
        RECT 4.000 112.900 295.600 114.900 ;
        RECT 4.000 112.860 296.000 112.900 ;
        RECT 4.000 110.860 295.600 112.860 ;
        RECT 4.000 110.820 296.000 110.860 ;
        RECT 4.000 110.140 295.600 110.820 ;
        RECT 4.400 108.820 295.600 110.140 ;
        RECT 4.400 108.780 296.000 108.820 ;
        RECT 4.400 108.140 295.600 108.780 ;
        RECT 4.000 106.780 295.600 108.140 ;
        RECT 4.000 106.740 296.000 106.780 ;
        RECT 4.000 104.740 295.600 106.740 ;
        RECT 4.000 104.700 296.000 104.740 ;
        RECT 4.000 102.700 295.600 104.700 ;
        RECT 4.000 102.660 296.000 102.700 ;
        RECT 4.000 100.660 295.600 102.660 ;
        RECT 4.000 99.940 296.000 100.660 ;
        RECT 4.000 98.580 295.600 99.940 ;
        RECT 4.400 97.940 295.600 98.580 ;
        RECT 4.400 97.900 296.000 97.940 ;
        RECT 4.400 96.580 295.600 97.900 ;
        RECT 4.000 95.900 295.600 96.580 ;
        RECT 4.000 95.860 296.000 95.900 ;
        RECT 4.000 93.860 295.600 95.860 ;
        RECT 4.000 93.820 296.000 93.860 ;
        RECT 4.000 91.820 295.600 93.820 ;
        RECT 4.000 91.780 296.000 91.820 ;
        RECT 4.000 89.780 295.600 91.780 ;
        RECT 4.000 89.740 296.000 89.780 ;
        RECT 4.000 87.740 295.600 89.740 ;
        RECT 4.000 87.700 296.000 87.740 ;
        RECT 4.000 87.020 295.600 87.700 ;
        RECT 4.400 85.700 295.600 87.020 ;
        RECT 4.400 85.660 296.000 85.700 ;
        RECT 4.400 85.020 295.600 85.660 ;
        RECT 4.000 83.660 295.600 85.020 ;
        RECT 4.000 83.620 296.000 83.660 ;
        RECT 4.000 81.620 295.600 83.620 ;
        RECT 4.000 81.580 296.000 81.620 ;
        RECT 4.000 79.580 295.600 81.580 ;
        RECT 4.000 79.540 296.000 79.580 ;
        RECT 4.000 77.540 295.600 79.540 ;
        RECT 4.000 77.500 296.000 77.540 ;
        RECT 4.000 75.500 295.600 77.500 ;
        RECT 4.000 75.460 296.000 75.500 ;
        RECT 4.400 74.780 296.000 75.460 ;
        RECT 4.400 73.460 295.600 74.780 ;
        RECT 4.000 72.780 295.600 73.460 ;
        RECT 4.000 72.740 296.000 72.780 ;
        RECT 4.000 70.740 295.600 72.740 ;
        RECT 4.000 70.700 296.000 70.740 ;
        RECT 4.000 68.700 295.600 70.700 ;
        RECT 4.000 68.660 296.000 68.700 ;
        RECT 4.000 66.660 295.600 68.660 ;
        RECT 4.000 66.620 296.000 66.660 ;
        RECT 4.000 64.620 295.600 66.620 ;
        RECT 4.000 64.580 296.000 64.620 ;
        RECT 4.000 63.900 295.600 64.580 ;
        RECT 4.400 62.580 295.600 63.900 ;
        RECT 4.400 62.540 296.000 62.580 ;
        RECT 4.400 61.900 295.600 62.540 ;
        RECT 4.000 60.540 295.600 61.900 ;
        RECT 4.000 60.500 296.000 60.540 ;
        RECT 4.000 58.500 295.600 60.500 ;
        RECT 4.000 58.460 296.000 58.500 ;
        RECT 4.000 56.460 295.600 58.460 ;
        RECT 4.000 56.420 296.000 56.460 ;
        RECT 4.000 54.420 295.600 56.420 ;
        RECT 4.000 54.380 296.000 54.420 ;
        RECT 4.000 52.380 295.600 54.380 ;
        RECT 4.000 52.340 296.000 52.380 ;
        RECT 4.400 50.340 295.600 52.340 ;
        RECT 4.000 49.620 296.000 50.340 ;
        RECT 4.000 47.620 295.600 49.620 ;
        RECT 4.000 47.580 296.000 47.620 ;
        RECT 4.000 45.580 295.600 47.580 ;
        RECT 4.000 45.540 296.000 45.580 ;
        RECT 4.000 43.540 295.600 45.540 ;
        RECT 4.000 43.500 296.000 43.540 ;
        RECT 4.000 41.500 295.600 43.500 ;
        RECT 4.000 41.460 296.000 41.500 ;
        RECT 4.000 40.780 295.600 41.460 ;
        RECT 4.400 39.460 295.600 40.780 ;
        RECT 4.400 39.420 296.000 39.460 ;
        RECT 4.400 38.780 295.600 39.420 ;
        RECT 4.000 37.420 295.600 38.780 ;
        RECT 4.000 37.380 296.000 37.420 ;
        RECT 4.000 35.380 295.600 37.380 ;
        RECT 4.000 35.340 296.000 35.380 ;
        RECT 4.000 33.340 295.600 35.340 ;
        RECT 4.000 33.300 296.000 33.340 ;
        RECT 4.000 31.300 295.600 33.300 ;
        RECT 4.000 31.260 296.000 31.300 ;
        RECT 4.000 29.260 295.600 31.260 ;
        RECT 4.000 29.220 296.000 29.260 ;
        RECT 4.400 27.220 295.600 29.220 ;
        RECT 4.000 27.180 296.000 27.220 ;
        RECT 4.000 25.180 295.600 27.180 ;
        RECT 4.000 24.460 296.000 25.180 ;
        RECT 4.000 22.460 295.600 24.460 ;
        RECT 4.000 22.420 296.000 22.460 ;
        RECT 4.000 20.420 295.600 22.420 ;
        RECT 4.000 20.380 296.000 20.420 ;
        RECT 4.000 18.380 295.600 20.380 ;
        RECT 4.000 18.340 296.000 18.380 ;
        RECT 4.000 17.660 295.600 18.340 ;
        RECT 4.400 16.340 295.600 17.660 ;
        RECT 4.400 16.300 296.000 16.340 ;
        RECT 4.400 15.660 295.600 16.300 ;
        RECT 4.000 14.300 295.600 15.660 ;
        RECT 4.000 14.260 296.000 14.300 ;
        RECT 4.000 12.260 295.600 14.260 ;
        RECT 4.000 12.220 296.000 12.260 ;
        RECT 4.000 10.220 295.600 12.220 ;
        RECT 4.000 10.180 296.000 10.220 ;
        RECT 4.000 8.180 295.600 10.180 ;
        RECT 4.000 8.140 296.000 8.180 ;
        RECT 4.000 6.780 295.600 8.140 ;
        RECT 4.400 6.140 295.600 6.780 ;
        RECT 4.400 6.100 296.000 6.140 ;
        RECT 4.400 4.780 295.600 6.100 ;
        RECT 4.000 4.100 295.600 4.780 ;
        RECT 4.000 4.060 296.000 4.100 ;
        RECT 4.000 2.895 295.600 4.060 ;
  END
END wrapped_bfloat16
END LIBRARY

